package proc_params is
end proc_params;
