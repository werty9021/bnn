package tta_core_params is
  constant fu_LSU1_addrw_g : integer := 14;
end tta_core_params;
