package tta0_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 30;
  constant fu_LSU_inp_dataw : integer := 32;
  constant fu_LSU_inp_addrw : integer := 24;
end tta0_params;
