package tta_core_toplevel_params is
  constant fu_LSU1_addrw_g : integer := 16;
  constant fu_DMA_addr_width_g : integer := 32;
  constant fu_DMA_data_width_g : integer := 32;
end tta_core_toplevel_params;
