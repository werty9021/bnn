package tta_core_toplevel_params is
  constant fu_DMA_addr_width_g : integer := 32;
  constant fu_DMA_data_width_g : integer := 32;
  constant fu_dmem_LSU_addrw_g : integer := 13;
end tta_core_toplevel_params;
