library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.tta0_imem_mau.all;

package tta0_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"0001011111110111111110111111111111101000010100000000000000011111100000000011000",
"0001011111110111111100000000010011111111111111100000000000000000100000000100100",
"0001011111110111111101000000110001011000001011000000000000000000000001111100000",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111100000000000000000000001010100000",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111100000000000000000010000000011001",
"0001011111110111111000000001010001000000101011000000000000000000000001011100001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111100000000010010000000010100000000000000000011100000000100100",
"0001011111110111111101000000110001011000010010000000000000000010111111100000000",
"0001011111110111111101000000101101000000010010000000000000000010100000000000000",
"0001011111110111111100000001000001111111111111100000000000000100110000000010011",
"0001011111110111111110111111111111111111111111100000000000000100111000000010011",
"0001011111110111111110111111111111111111111111100000000000000101000000000010011",
"0001011111110111111110111111111111111111111111100000000000000101001000000010011",
"0001011111110011100101000000101111111111111111100000000000000010000000000000000",
"0001011111110011100101000000101111000000010010000000000000000001100000000000000",
"0001011111110011100101000000101111000000010010000000000000000001000000000000000",
"0001011111110011100101000000101111000000010010000000000000000000100000000000000",
"0001011111110111111110111111111111111111111111100000000000000101010000000010000",
"0001011111110111111110111111111111111111111111100000000000000101100000000010000",
"0001011111110111111110111111111111111111111111100000000000000000000100000100001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001001110010111111101000000101001111111111111111101111111111111111111111111111",
"0001001110010111111100000000101001000000010010000000000000000010100000000000000",
"0001011111110111111101000000100111000000010010000000000000000010000000000000000",
"0001011111110111111101000000100111111111111111100000000000000000100000000011001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110011000110111111111111111111111111111101111111111111111111111111111",
"0001011111110000101110111111111111111111111111111101111111111111111111111111111",
"0001011111111011100100000010101111111111111111111101111111111111111111111111111",
"0001011111110111111100000001000000000000101100100000000000000010100000000000000",
"0001011111110111111101000000100111000000010010000000000000000001000000000011100",
"0001011111110111111110111111111111111111111111100000000000000000000000001101100",
"0001011111110111111110111111111111111111111111100000000000000000100000000000000",
"0001011111110111111101000000100001111111111111111101111111111111111111111111111",
"0001011111110000110110111111111111111111111111111101111111111111111111111111111",
"0001011111111011100100001000101111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111100000100000000000000000001101100",
"0001000011110111111110111111111111111111111111111101111111111111111111111111111",
"0001101110010111111110111111111111111111111111100000000000000001100000000010100",
"0001011111110111111100000001000001111111111111100000000000000000100000000000000",
"0001011111110111111101000000100001111111111111100000000000000010000000000011001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001000100010111111110111111111111111111111111111101111111111111111111111111111",
"0001101110010111111100000010101111111111111111111101111111111111111111111111111",
"0001011111110111111100000001000001111111111111100000000000000010100000000000000",
"0001011111110111111101000000100111111111111111100000000000000000000110110101100",
"0001011111110111111110111111111111111111111111100000000000000000000000000101000",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110000010110111111111111111111111111111101111111111111111111111111111",
"0001011111111011100110111111111111111111111111100000000000000010100000000010111",
"0001011111110111111100000000100001111111111111100000000000000000000111010101100",
"0001011111110111111110111111111111111111111111100000000000000000000000000101000",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001000001110111111110111111111111111111111111111101111111111111111111111111111",
"0001101110010111111110111111111111111111111111100000000000000010100000000010111",
"1001011111110111111100000001000000000000010100011111111111111111111111111111100",
"1001011111110111111100100000000001111111111111111111111111111111111111111111100",
"0001011111110111111101000000101101000000010010000000000000000001100000000000000",
"0001011111110111111101000000100111000000010010000000000000000001000000000000000",
"0001011111110111111101000000100111001000000000000000100000000000000000000100100",
"1001011111110111111101000000111001000000010010011111111111111111111111111111100",
"0001011111110111111100100000000001111111111111111101111111111111111111111111111",
"0001011111110010000110111111111111111111111111111101111111111111111111111111111",
"0001011111110010100110111111111111111111111111111101111111111111111111111111111",
"0001011111100000001110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111101100001010001000010001011000000000000000011000000000011100",
"0001011111110111111101000000100101111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001010001000010001011011101111111111111111111111111111",
"1001011111110111111100000001000000000000010100011111111111111111111111111111000",
"1001011111110111111100100000000001111111111111111111111111111111111111111111000",
"0001011111110111111101000000101101000000010010000000000000000001000000000000000",
"0001011111110111111101000000100111000000010010000000000000000001100000000000000",
"0001011111110111111101000000100111001000000000000000100000000000000000000100100",
"1001011111110111111101000000111001000000010010011111111111111111111111111111000",
"0001011111110111111100100000000001111111111111111101111111111111111111111111111",
"0001011111110010000110111111111111111111111111111101111111111111111111111111111",
"0001011111110010100110111111111111111111111111111101111111111111111111111111111",
"0001011111100000001110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111101100001010001000010001011000000000000000011100000000011100",
"0001011111110111111101000000100101111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001010001000010001011011101111111111111111111111111111",
"1001011111110111111100000001000000000000010100011111111111111111111111111110100",
"1001011111110111111100100000000001000000001000011111111111111111111111111110100",
"0001011111110111111101000000101101000000010010000000000000000000100000000000000",
"0001011111110111111101000000100001001000000000000000100000000000000000000100100",
"1001011111110111111101000000111001000000010010011111111111111111111111111110100",
"0001001000110111111100100000000001111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001001100010111111110111111111111111111111111111101111111111111111111111111111",
"0000010000010111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111101100001010001000010001011000000000000000011100000100011100",
"0001011111110111111101000000100101111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001010001000010001011011101111111111111111111111111111",
"1001011111110111111100000001000000000000010100011111111111111111111111111110000",
"1001011111110111111100100000000001000000001000011111111111111111111111111110000",
"0001011111110111111101000000101101000000010010000000000000000000100000000000000",
"0001011111110111111101000000100001001000000000000000100000000000000000000100100",
"1001011111110111111101000000111001000000010010011111111111111111111111111110000",
"0001001100010111111100100000000001111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001000000010111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111101100001010001000010001011000000000000000011100001000011100",
"0001011111110111111101000000100101111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001010001000010001011011101111111111111111111111111111",
"0001011111110111111110111111111111111111111111100000000000000000010001010100001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111100000001000001111111111111100000000000000010100000000000000",
"0001011111110111111101000000100111000000010010000000000000000010000000000000000",
"0001011111110111111101000000100111000000010010000000000000000000100000000000000",
"0001011111110111111101000000100001111111111111100000000000000100000000000011001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110010000110111111111111111111111111111101111111111111111111111111111",
"0001011111110010100110111111111111111111111111111101111111111111111111111111111",
"0001001100000000100110111111111111111111111111111101111111111111111111111111111",
"0001101110010111111100000010101001111111111111111101111111111111111111111111111",
"1001011111110111111100000001000000000000010100011111111111111111111111111101100",
"1001011111110111111100100000000001111111111111111111111111111111111111111101100",
"0001011111110111111101000000101101000000010010000000000000000000100000000000000",
"0001011111110111111101000000100001001000000000000000100000000000000000000100100",
"1001011111110111111101000000111001000000010010011111111111111111111111111101100",
"0001011111110111111100100000000001111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001000100110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111101100001010001000010001011000000000000000100010000000011100",
"0001011111110111111101000000100101111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001010001000010001011011101111111111111111111111111111",
"0001011111110111111100000001000001000000001000000000000000000000100000000000000",
"0001011111110111111101000000100001000000010010000000000000000010100000000000000",
"0001011111110111111101000000100111111111111111100000000000000100100000000011001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001001000110111111110111111111111111111111111111101111111111111111111111111111",
"0001001000010111111110111111111111111111111111111101111111111111111111111111111",
"0000001010010011000110111111111111111111111111111101111111111111111111111111111",
"0000010101010111111110111111111111111111111111111101111111111111111111111111111",
"0001101110011010000100000010101111111111111111111101111111111111111111111111111",
"0001011111110111111100000001000001101000001111100000000000000100101000000010010",
"0001011111110111111110111111111111111111111111100000000000000011100000000000000",
"0001011111110111111101000000110001111111111111111101111111111111111111111111111",
"0001011111110111111110111111111111111111111111100000100000000000000000111100001",
"0001011111110111111110111111111111111111111111111101111111111111111111111111111",
"0001011111110111111110000001000000000000100000011101111111111111111111111111111",
"0001011111110111111101000000110011011000010100000000000000000100101000100010110");

end tta0_imem_image;
