package tta_core_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 82;
end tta_core_imem_mau;
